MODULE aktuell
 
TITLE 'Abelprojekt'
 
@dcset
 
DECLARATIONS
"Eingänge"
G0,G1,G2,G3,takt,Motorstart PIN 91,93,94,98,88,17;
M0,M1,M2,M3 PIN 31,30,29,28;
 
"Ausgänge"
Q0 PIN 56 ISTYPE 'BUFFER,REG';
Q1 PIN 55 istype 'BUFFER,REG';
Q2 PIN 54 istype 'BUFFER,REG';
Q3 PIN 53 istype 'Buffer,REG';
aa,bb,cc,dd,ee,ff,gg PIN 81,79,80,85,87,84,86 istype 'Buffer,COM';
a,b,c,d,e,f,g PIN 67,65,66,70,72,69,71 ISTYPE 'BUFFER,COM';
AnMotor,DrehRichtung  PIN 37,36 ISTYPE 'BUFFER,COM';
 
 
C3 NODE ISTYPE 'BUFFER,COM';
T0,T1,T2,T3,T4 node ISTYPE 'BUFFER,COM';
 
x =.X.;
 
 
"Set"
Zustandreg = [Q3,Q2,Q1,Q0];
Bin = [Q3,Q2,Q1,Q0];
Gray = [G3,G2,G1,G0];
Maus = [M3,M2,M1,M0];
bcd = [T0,T1,T2,T3,T4];
IDLE =0;
Drive =1;
"gleich = (Bin != Maus);"
 
EQUATIONS
Zustandreg.CLK = takt;
"AnMotor = Motorstart;"
when Bin != Maus then AnMotor = 1;
 
"State_DIAGRAM Zustandreg;"
"state IDLE: "
"If Bin != Maus then AnMotor else IDLE;"
"state Drive:"
"AnMotor =1; "
"goto IDLE;"
 
 
Truth_Table (Gray -> Bin)
[0,0,0,0]->[0,0,0,0];
[0,0,0,1]->[0,0,0,1];
[0,0,1,1]->[0,0,1,0];
[0,0,1,0]->[0,0,1,1];
[0,1,1,0]->[0,1,0,0];
[0,1,1,1]->[0,1,0,1];
[0,1,0,1]->[0,1,1,0];
[0,1,0,0]->[0,1,1,1];
[1,1,0,0]->[1,0,0,0];
[1,1,0,1]->[1,0,0,1];
[1,1,1,1]->[1,0,1,0];
[1,1,1,0]->[1,0,1,1];
[1,0,1,0]->[1,1,0,0];
[1,0,1,1]->[1,1,0,1];
[1,0,0,1]->[1,1,1,0];
[1,0,0,0]->[1,1,1,1];
 
Truth_Table (Bin -> bcd)
[0,0,0,0]->[0,0,0,0,0];
[0,0,0,1]->[0,0,0,0,1];
[0,0,1,0]->[0,0,0,1,0];
[0,0,1,1]->[0,0,0,1,1];
[0,1,0,0]->[0,0,1,0,0];
[0,1,0,1]->[0,0,1,0,1];
[0,1,1,0]->[0,0,1,1,0];
[0,1,1,1]->[0,0,1,1,1];
[1,0,0,0]->[0,1,0,0,0];
[1,0,0,1]->[0,1,0,0,1];
[1,0,1,0]->[1,0,0,0,0];
[1,0,1,1]->[1,0,0,0,1];
[1,1,0,0]->[1,0,0,1,0];
[1,1,0,1]->[1,0,0,1,1];
[1,1,1,0]->[1,0,1,0,0];
[1,1,1,1]->[1,0,1,0,1];
 
TRUTH_TABLE (bcd ->[a,b,c,d,e,f,g])  "BCD -> 7 Segment"
[0,0,0,0,0]->[1,1,1,1,1,1,0];
[0,0,0,0,1]->[0,1,1,0,0,0,0];
[0,0,0,1,0]->[1,1,0,1,1,0,1];
[0,0,0,1,1]->[1,1,1,1,0,0,1];
[0,0,1,0,0]->[0,1,1,0,0,1,1];
[0,0,1,0,1]->[1,0,1,1,0,1,1];
[0,0,1,1,0]->[1,0,1,1,1,1,1];
[0,0,1,1,1]->[1,1,1,0,0,0,0];
[0,1,0,0,0]->[1,1,1,1,1,1,1];
[0,1,0,0,1]->[1,1,1,1,1,0,1];
[1,0,0,0,0]->[1,1,1,1,1,1,0];
[1,0,0,0,1]->[0,1,1,0,0,0,0];
[1,0,0,1,0]->[1,1,0,1,1,0,1];
[1,0,0,1,1]->[1,1,1,1,0,0,1];
[1,0,1,0,0]->[0,1,1,0,0,1,1];
[1,0,1,0,1]->[1,0,1,1,0,1,1];
 
TRUTH_TABLE (bcd ->[aa,bb,cc,dd,ee,ff,gg])  "BCD -> 7 Segment"
[0,0,0,0,0]->[0,0,0,0,0,0,0];
[0,0,0,0,1]->[0,0,0,0,0,0,0];
[0,0,0,1,0]->[0,0,0,0,0,0,0];
[0,0,0,1,1]->[0,0,0,0,0,0,0];
[0,0,1,0,0]->[0,0,0,0,0,0,0];
[0,0,1,0,1]->[0,0,0,0,0,0,0];
[0,0,1,1,0]->[0,0,0,0,0,0,0];
[0,0,1,1,1]->[0,0,0,0,0,0,0];
[0,1,0,0,0]->[0,0,0,0,0,0,0];
[0,1,0,0,1]->[0,0,0,0,0,0,0];
[1,0,0,0,0]->[0,1,1,0,0,0,0];
[1,0,0,0,1]->[0,1,1,0,0,0,0];
[1,0,0,1,0]->[0,1,1,0,0,0,0];
[1,0,0,1,1]->[0,1,1,0,0,0,0];
[1,0,1,0,0]->[0,1,1,0,0,0,0];
[1,0,1,0,1]->[0,1,1,0,0,0,0];
 
 
END