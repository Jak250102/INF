Module Test
 
Title 'Kreuz und Quer'
 
@dcset
 
Declarations

"Eingänge

Start, V_R, takt Pin 30,31,88;
 
"Ausgänge

Flip0,Flip1,Flip2,Flip3 pin 56,55,54,53 istype 'buffer.Reg';

a,b,c,d,e,f,g Pin 67,65,66,70,72,69,71 istype 'Buffer.com';
 
"Set

ff = [Flip3,Flip2,Flip1,Flip0];
 
equations

ff.clk = takt;

Truth_table ([Start,V_R,Flip3,Flip2,Flip1,Flip0] :> ff)

[0,0,0,0,0,0]:>[0,0,0,0];

[0,0,0,0,0,1]:>[0,0,0,1];

[0,0,0,0,1,0]:>[0,0,1,0];

[0,0,0,0,1,1]:>[0,0,1,1];

[0,0,0,1,0,0]:>[0,1,0,0];

[0,0,0,1,0,1]:>[0,1,0,1];

[0,0,0,1,1,0]:>[0,1,1,0];

[0,0,0,1,1,1]:>[0,1,1,1];

[0,0,1,0,0,0]:>[1,0,0,0];

[0,0,1,0,0,1]:>[1,0,0,1];

[0,1,0,0,0,0]:>[0,0,0,0];

[0,1,0,0,0,1]:>[0,0,0,1];

[0,1,0,0,1,0]:>[0,0,1,0];

[0,1,0,0,1,1]:>[0,0,1,1];

[0,1,0,1,0,0]:>[0,1,0,0];

[0,1,0,1,0,1]:>[0,1,0,1];

[0,1,0,1,1,0]:>[0,1,1,0];

[0,1,0,1,1,1]:>[0,1,1,1];

[0,1,1,0,0,0]:>[1,0,0,0];

[0,1,1,0,0,1]:>[1,0,0,1];

[1,0,0,0,0,0]:>[0,1,1,0];

[1,0,0,0,0,1]:>[0,1,0,0];

[1,0,0,0,1,0]:>[0,1,1,1];

[1,0,0,0,1,1]:>[0,0,0,0];

[1,0,0,1,0,0]:>[1,0,0,1];

[1,0,0,1,0,1]:>[1,0,0,0];

[1,0,0,1,1,0]:>[0,0,1,0];

[1,0,0,1,1,1]:>[0,0,0,1];

[1,0,1,0,0,0]:>[0,0,1,1];

[1,0,1,0,0,1]:>[0,1,0,1];

[1,1,0,0,0,0]:>[0,0,1,1];

[1,1,0,0,0,1]:>[0,1,1,1];

[1,1,0,0,1,0]:>[0,1,1,0];

[1,1,0,0,1,1]:>[1,0,0,0];

[1,1,0,1,0,0]:>[0,0,0,1];

[1,1,0,1,0,1]:>[1,0,0,1];

[1,1,0,1,1,0]:>[0,0,0,0];

[1,1,0,1,1,1]:>[0,0,1,0];

[1,1,1,0,0,0]:>[0,1,0,1];

[1,1,1,0,0,1]:>[0,1,0,0];
 
truth_table (ff -> [a,b,c,d,e,f,g])

0 -> [1,1,1,1,1,1,0];

1 -> [0,1,1,0,0,0,0];

2 -> [1,1,0,1,1,0,1];

3 -> [1,1,1,1,0,0,1];

4 -> [0,1,1,0,0,1,1];

5 -> [1,0,1,1,0,1,1];

6 -> [1,0,1,1,1,1,1];

7 -> [1,1,1,0,0,0,0];

8 -> [1,1,1,1,1,1,1];

9 -> [1,1,1,1,1,0,1];
 
 
end
 