MODULE test

TITLE 'test'
@dcset

DECLARATIONS

"Eingänge"
C0, C1, C2, C3 Pin 31, 30, 29, 28;

tmp1, tmp2, tmp3 NODE ISTYPE 'BUFFER,COM';

"Ausgänge"
J, Y, Z, U, V, W, S Pin 81, 79, 80, 85, 87, 84, 86 ISTYPE 'BUFFER,COM';
x=.X.;
"Set"
set1=[C3, C2, C1, C0];

"Equations" "enteweder Equations oder Truth Table"
"Peter = !C0;"

"TRUTH_TABLE ([C3, C2, C1, C0] -> [J, Y, Z, U, V, W, S])"
"[0, 0, 0, 0] -> [1, 1, 1, 1, 1, 1, 0];"
"[0, 0, 0, 1] -> [0, 1, 1, 0, 0, 0, 0];"
"[0, 0, 1, 0] -> [1, 1, 0, 1, 1, 0, 1];"
"[0, 0, 1, 1] -> [1, 1, 1, 1, 0, 0, 1];"
"[0, 1, 0, 0] -> [0, 1, 1, 0, 0, 1, 1];"
"[0, 1, 0, 1] -> [1, 0, 1, 1, 0, 1, 1];"
"[0, 1, 1, 0] -> [1, 0, 1, 1, 1, 1, 1];"
"[0, 1, 1, 1] -> [1, 1, 1, 0, 0, 0, 0];"
"[1, 0, 0, 0] -> [1, 1, 1, 1, 1, 1, 1];"
"[1, 0, 0, 1] -> [1, 1, 1, 1, 0, 1, 1];"
"[1, 0, 1, 0] -> [1, 1, 0, 1, 1, 1, 1];"
"[1, 0, 1, 1] -> [1, 1, 1, 1, 0, 1, 1];"
"[1, 1, 0, 0] -> [1, 1, 1, 1, 0, 1, 1];"
"[1, 1, 0, 1] -> [1, 0, 1, 1, 0, 1, 1];"
"[1, 1, 1, 0] -> [1, 0, 1, 1, 1, 1, 1];"
"[1, 1, 1, 1] -> [1, 1, 1, 1, 0, 1, 1];"

TRUTH_TABLE (set1 -> [J, Y, Z, U, V, W, S])
0 -> [1, 1, 1, 1, 1, 1, 0];
1 -> [0, 1, 1, 0, 0, 0, 0];
2 -> [1, 1, 0, 1, 1, 0, 1];
3 -> [1, 1, 1, 1, 0, 0, 1];
4 -> [0, 1, 1, 0, 0, 1, 1];
5 -> [1, 0, 1, 1, 0, 1, 1];
6 -> [1, 0, 1, 1, 1, 1, 1];
7 -> [1, 1, 1, 0, 0, 0, 0];
8 -> [1, 1, 1, 1, 1, 1, 1];
9 -> [1, 1, 1, 1, 0, 1, 1];
10 -> [1, 1, 0, 1, 1, 1, 1];
11 -> [1, 1, 1, 1, 0, 1, 1];
12 -> [1, 1, 1, 1, 0, 1, 1];
13 -> [1, 0, 1, 1, 0, 1, 1];
14 -> [1, 0, 1, 1, 1, 1, 1];
15 -> [1, 1, 1, 1, 0, 1, 1];

END