MODULE aktuell

TITLE 'aktuell'


@dcset

DECLARATIONS
takt PIN 88; 

ff1,ff2,ff3 PIN 61,60,59 ISTYPE 'BUFFER, REG';

ff = [ff1,ff2,ff3];" SET

EQUATIONS
ff.clk = takt; "Takt auf alle ffs im SET legen 

TRUTH_TABLE

(ff :> ff)
0 :> 4;
1 :> 0;
2 :> 6;
3 :> 7;
4 :> 2;
5 :> 3;
6 :> 5;
7 :> 1;

TRUTH_TABLE
(ff ->[a,b,c,d,e,f,g]);
[0,0,0,0]->[1,1,1,1,1,1,0];
[0,0,0,1]->[0,1,1,0,0,0,0];
[0,0,1,0]->[1,1,0,1,1,0,1];
[0,0,1,1]->[1,1,1,1,0,0,1];
[0,1,0,0]->[0,1,1,0,0,1,1];
[0,1,0,1]->[1,0,1,1,0,1,1];
[0,1,1,0]->[1,0,1,1,1,1,1];
[0,1,1,1]->[1,1,1,0,0,0,0];
[1,0,0,0]->[1,1,1,1,1,1,1];
[1,0,0,1]->[1,1,1,1,0,1,1];
[1,0,1,0]->[x,x,x,x,x,x,x];
[1,0,1,1]->[x,x,x,x,x,x,x];
[1,1,0,0]->[x,x,x,x,x,x,x];
[1,1,0,1]->[x,x,x,x,x,x,x];
[1,1,1,0]->[x,x,x,x,x,x,x];
[1,1,1,1]->[x,x,x,x,x,x,x];


END
