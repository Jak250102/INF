MODULE aktuell

TITLE 'aktuell'


@dcset

DECLARATIONS
takt PIN 88; 
S1,S2 PIN 30,31;
A, B, C, D, E, F, G Pin 81, 79, 80, 85, 87, 84, 86 ISTYPE 'BUFFER,COM';

ff1,ff2,ff3,ff4 PIN ISTYPE 'BUFFER, REG';

ff = [ff1,ff2,ff3,ff4];" SET"

EQUATIONS
ff.clk = takt; "Takt auf alle ffs im SET legen "

TRUTH_TABLE

([S1,S2,ff1,ff2,ff3,ff4] :> ff ) " Vor dem Takt :> Nach dem Takt"
"---------------
" vorwaerts 
[0,0,0,0,0,0] :> 1;
[0,0,0,0,0,1] :> 2;
[0,0,0,0,1,0] :> 3;
[0,0,0,0,1,1] :> 4;
[0,0,0,1,0,0] :> 5;
[0,0,0,1,0,1] :> 6;
[0,0,0,1,1,0] :> 7;
[0,0,0,1,1,1] :> 8;
[0,0,1,0,0,0] :> 9;
[0,0,1,0,0,1] :> 0;

"---------------"


" Zaehler stoppt"
[1,0,0,0,0,0] :> 0;
[1,0,0,0,0,1] :> 1;
[1,0,0,0,1,0] :> 2;
[1,0,0,0,1,1] :> 3;
[1,0,0,1,0,0] :> 4;
[1,0,0,1,0,1] :> 5;
[1,0,0,1,1,0] :> 6;
[1,0,0,1,1,1] :> 7;
[1,0,1,0,0,0] :> 8;
[1,0,1,0,0,1] :> 9;
"---------------"
"Rueckwaerts"
[0,1,0,0,0,0] :> 9;
[0,1,0,0,0,1] :> 0;
[0,1,0,0,1,0] :> 1;
[0,1,0,0,1,1] :> 2;
[0,1,0,1,0,0] :> 3;
[0,1,0,1,0,1] :> 4;
[0,1,0,1,1,0] :> 5;
[0,1,0,1,1,1] :> 6;
[0,1,1,0,0,0] :> 7;
[0,1,1,0,0,1] :> 8;
[0,1,1,0,1,0] :> 9;



TRUTH_TABLE (ff -> [A, B, C, D, E, F, G])
  0 -> [1, 1, 1, 1, 1, 1, 0];
  1 -> [0, 1, 1, 0, 0, 0, 0];
  2 -> [1, 1, 0, 1, 1, 0, 1];
  3 -> [1, 1, 1, 1, 0, 0, 1];
  4 -> [0, 1, 1, 0, 0, 1, 1];
  5 -> [1, 0, 1, 1, 0, 1, 1];
  6 -> [1, 0, 1, 1, 1, 1, 1];
  7 -> [1, 1, 1, 0, 0, 0, 0];
  8 -> [1, 1, 1, 1, 1, 1, 1];
  9 -> [1, 1, 1, 1, 0, 1, 1];
  



END
